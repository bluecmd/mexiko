//////////////////////////////////////////////////////////////////////
//
// Xilinx specific 10G Ethernet PHY module
// Logic shared between 4 lanes in one bank. Based on the example design.
//
// Copyright (C) 2014 Christian Svensson <blue@cmd.nu>
//
//////////////////////////////////////////////////////////////////////
//
// This source file may be used and distributed without
// restriction provided that this copyright statement is not
// removed from the file and that any derivative work contains
// the original copyright notice and the associated disclaimer.
//
// This source file is free software; you can redistribute it
// and/or modify it under the terms of the GNU Lesser General
// Public License as published by the Free Software Foundation;
// either version 3 of the License, or (at your option) any
// later version.
//
// This source is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied
// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
// PURPOSE.  See the GNU Lesser General Public License for more
// details.
//
// You should have received a copy of the GNU Lesser General
// Public License along with this source; if not, download it
// from http://www.opencores.org/lgpl.shtml
//
//////////////////////////////////////////////////////////////////////

module  xilinx_phy10g_quad_logic (
  input  refclk_i,
  input  qpllreset_i,
  output qplllock_o,
  output qplloutclk_o,
  output qplloutrefclk_o
);
  localparam QPLL_FBDIV_TOP =  66;

  localparam QPLL_FBDIV_IN  =  (QPLL_FBDIV_TOP == 16)  ? 10'b0000100000 :
    (QPLL_FBDIV_TOP == 20)  ? 10'b0000110000 :
    (QPLL_FBDIV_TOP == 32)  ? 10'b0001100000 :
    (QPLL_FBDIV_TOP == 40)  ? 10'b0010000000 :
    (QPLL_FBDIV_TOP == 64)  ? 10'b0011100000 :
    (QPLL_FBDIV_TOP == 66)  ? 10'b0101000000 :
    (QPLL_FBDIV_TOP == 80)  ? 10'b0100100000 :
    (QPLL_FBDIV_TOP == 100) ? 10'b0101110000 : 10'b0000000000;

  localparam QPLL_FBDIV_RATIO = (QPLL_FBDIV_TOP == 16)  ? 1'b1 :
    (QPLL_FBDIV_TOP == 20)  ? 1'b1 :
    (QPLL_FBDIV_TOP == 32)  ? 1'b1 :
    (QPLL_FBDIV_TOP == 40)  ? 1'b1 :
    (QPLL_FBDIV_TOP == 64)  ? 1'b1 :
    (QPLL_FBDIV_TOP == 66)  ? 1'b0 :
    (QPLL_FBDIV_TOP == 80)  ? 1'b1 :
    (QPLL_FBDIV_TOP == 100) ? 1'b1 : 1'b1;

  wire            tied_to_ground_i;
  wire    [63:0]  tied_to_ground_vec_i;
  wire            tied_to_vcc_i;
  wire    [63:0]  tied_to_vcc_vec_i;

  assign tied_to_ground_i             = 1'b0;
  assign tied_to_ground_vec_i         = 64'h0000000000000000;
  assign tied_to_vcc_i                = 1'b1;
  assign tied_to_vcc_vec_i            = 64'hffffffffffffffff;

  wire gt0_gtrefclk0_common_in;
  wire gt0_qpllreset_in;
  wire gt0_qplllock_out;
  wire gt0_qplloutclk_i;
  wire gt0_qplloutrefclk_i;

  assign gt0_gtrefclk0_common_in = refclk_i;
  assign gt0_qpllreset_in = qpllreset_i;
  assign qplllock_o = gt0_qplllock_out;
  assign qplloutclk_o = gt0_qplloutclk_i;
  assign qplloutrefclk_o = gt0_qplloutrefclk_i;

  GTXE2_COMMON # (
    /* Simulation attributes */
    .SIM_RESET_SPEEDUP   ("false"),
    .SIM_QPLLREFCLK_SEL  (3'b001),
    .SIM_VERSION         ("4.0"),
    /* COMMON BLOCK Attributes */
    .BIAS_CFG                               (64'h0000040000001000),
    .COMMON_CFG                             (32'h00000000),
    .QPLL_CFG                               (27'h0680181),
    .QPLL_CLKOUT_CFG                        (4'b0000),
    .QPLL_COARSE_FREQ_OVRD                  (6'b010000),
    .QPLL_COARSE_FREQ_OVRD_EN               (1'b0),
    .QPLL_CP                                (10'b0000011111),
    .QPLL_CP_MONITOR_EN                     (1'b0),
    .QPLL_DMONITOR_SEL                      (1'b0),
    .QPLL_FBDIV                             (QPLL_FBDIV_IN),
    .QPLL_FBDIV_MONITOR_EN                  (1'b0),
    .QPLL_FBDIV_RATIO                       (QPLL_FBDIV_RATIO),
    .QPLL_INIT_CFG                          (24'h000006),
    .QPLL_LOCK_CFG                          (16'h21E8),
    .QPLL_LPF                               (4'b1111),
    .QPLL_REFCLK_DIV                        (1)
  ) gtxe2_common_i (
    /* Common Block - Dynamic Reconfiguration Port (DRP) */
    .DRPADDR                        (tied_to_ground_vec_i[7:0]),
    .DRPCLK                         (tied_to_ground_i),
    .DRPDI                          (tied_to_ground_vec_i[15:0]),
    .DRPDO                          (),
    .DRPEN                          (tied_to_ground_i),
    .DRPRDY                         (),
    .DRPWE                          (tied_to_ground_i),
    /* Common Block - Ref Clock Ports */
    .GTGREFCLK                      (tied_to_ground_i),
    .GTNORTHREFCLK0                 (tied_to_ground_i),
    .GTNORTHREFCLK1                 (tied_to_ground_i),
    .GTREFCLK0                      (gt0_gtrefclk0_common_in),
    .GTREFCLK1                      (tied_to_ground_i),
    .GTSOUTHREFCLK0                 (tied_to_ground_i),
    .GTSOUTHREFCLK1                 (tied_to_ground_i),
    /* Common Block - Clocking Ports */
    .QPLLOUTCLK                     (gt0_qplloutclk_i),
    .QPLLOUTREFCLK                  (gt0_qplloutrefclk_i),
    .REFCLKOUTMONITOR               (),
    /* Common Block - QPLL Ports */
    .QPLLDMONITOR                   (),
    .QPLLFBCLKLOST                  (),
    .QPLLLOCK                       (gt0_qplllock_out),
    .QPLLLOCKDETCLK                 (1'b0),
    .QPLLLOCKEN                     (tied_to_vcc_i),
    .QPLLOUTRESET                   (tied_to_ground_i),
    .QPLLPD                         (tied_to_ground_i),
    .QPLLREFCLKLOST                 (),
    .QPLLREFCLKSEL                  (3'b001),
    .QPLLRESET                      (gt0_qpllreset_in),
    .QPLLRSVD1                      (16'b0000000000000000),
    .QPLLRSVD2                      (5'b11111),
    /* QPLL Ports */
    .BGBYPASSB                      (tied_to_vcc_i),
    .BGMONITORENB                   (tied_to_vcc_i),
    .BGPDB                          (tied_to_vcc_i),
    .BGRCALOVRD                     (5'b00000),
    .PMARSVD                        (8'b00000000),
    .RCALENB                        (tied_to_vcc_i)
  );
endmodule
