`define USE_EMERGENCY_CLK