`define MOR1KX